/*
 * A Testbench of the Wrapper for BCH Encoder
 *
 * Copyright 2015 - Lix Wei <ultracold273@outlook.com>
 * Encoder Module comes from Russ Dill
 *
 * Encodes the bits and save the ecc bits to outside memory
 */

`include "../bch_verilog/bch_params.vh"
`include "../bch_verilog/bch_defs.vh"

module test_bch_wrapper_encode();
localparam 
bch_wrapper_encoder #() (
);
endmodule
